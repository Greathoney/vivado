module bin2seg(
input	wire	[3:0]	bin,

output	reg		[7:0]	seg
);

always @(bin)
begin
	case(bin)
		////////////////////////////////////////////
		//
		//
		//
		//
		// Coding here!
		//
		//
		//
		//
		//
		////////////////////////////////////////////
	endcase
end

endmodule
